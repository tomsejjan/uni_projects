--! \file testbench.vhdl
--! \brief Definice entity a architektury Testbench urcene pro testovani DUT (Device Under Test) komponent: Led7seg_adder3, Adder3, Led7seg_decoder_hex

--! Zavedena standardni knihovna \c IEEE
LIBRARY ieee;
--! Zpristupnen balik \c std_logic_1164 z knihovny \c IEEE pro podporu 9-ti stavove logiky
USE ieee.std_logic_1164.ALL;
--! Zpristupnen balik \c numeric_std z knihovny \c IEEE pro podporu konverze cisel dle IEEE 1076.3
USE ieee.numeric_std.ALL;

--LIBRARY work;
--! Zpristupnen cely balik \c pkg_bpc_los z pracovni knihovny \c work pro podporu zobrazeni stavu 7-seg displeje
USE work.pkg_bpc_los.ALL;

--! \brief Definice entity Testbench
--! \details Entita Testbench overuje spravnost komponent: Led7seg_adder3, Adder3, Led7seg_decoder_hex.
ENTITY Testbench IS
	-- Entita Testbench nebude mit zadne vstupy ani vystupy
END Testbench;

--! \brief Definice architektury entity Testbench
--! \details Architektura entity Testbench overuje spravnost komponent: Led7seg_adder3, Adder3, Led7seg_decoder_hex.
ARCHITECTURE Behavioral of Testbench IS

	CONSTANT stimulus_step_c: delay_length := 10 ns;	--! Definice a inicializace konstanty simulace

	--! \brief DUT (Device Under Test) komponenta Led7seg_adder3
	COMPONENT Led7seg_adder3 IS
		PORT(
			a:   in std_logic_vector(2 downto 0);		-- Deklarace vstupu: a[2:0]
			b:   in std_logic_vector(2 downto 0);		-- Deklarace vstupu: b[2:0]
			cin: in std_logic;				-- Deklarace vstupu: carry in
			an:  out std_logic_vector(3 downto 0);		-- Deklarace vystupu: an[3:0]
			seg: out std_logic_vector(6 downto 0)		-- Deklarace vystupu: seg[6:0]
			);
	END COMPONENT Led7seg_adder3;

	SIGNAL a_in, b_in: std_logic_vector(2 DOWNTO 0) := (OTHERS => '0'); --! Definice signalu pripojenych na vstupy testovane komponenty
	SIGNAL c_in: std_logic := '0';					--! Definice signalu pripojeneho na vstupy testovane komponenty
	SIGNAL an_out: std_logic_vector(3 DOWNTO 0);	--! Definice signalu pripojenych na vystupy testovane komponenty (anody)
	SIGNAL seg_out: std_logic_vector(6 DOWNTO 0);	--! Definice signalu pripojenych na vystupy testovane komponenty (katody)

	-- Mapping alias to the internal signal and port with VHDL-2008 External name feature
	ALIAS dut_sum_result IS							--! Pripojeni na vnitrni signal \p sum_result_i testovane komponenty Led7seg_adder3
		<< SIGNAL .Testbench.dut.sum_result_i: std_logic_vector(3 DOWNTO 0) >>;
BEGIN
	-- Pripojime DUT komponentu Led7seg_adder3 na jednotlive stimuly pomoci jmenne asociace
	dut: Led7seg_adder3
		PORT MAP(
			a   => a_in,
			b   => b_in,
			cin => c_in,
			an  => an_out,
			seg => seg_out
			);

	--! \vhdlflow testbench_proc
	--! \test **Test #0 - #3**\n
	--!   Testujeme spravnou funkci Testujeme Adder3 a Led7seg_decoder_hex na prikladech (1+1+1, 4+2+0, 7+7+1)\n
	--! \test **Test #4 - #132**\n
	--!   Testujeme spravnou funkci Adder3 na vsech moznych kombinacich vstupu: a, b, cin.
	testbench_proc: PROCESS
	BEGIN
		REPORT "Test start." SEVERITY note;

		-- Testujeme Adder3 a Led7seg_decoder_hex
		REPORT "Testing Led7seg_adder3..." SEVERITY note;
		REPORT "1 + 1 + 1 =" SEVERITY note;
		a_in <= O"1";
		b_in <= O"1";
		c_in <= '1';
		WAIT FOR stimulus_step_c;
		led7seg_show_big(an_out, seg_out);

		REPORT "4 + 2 + 0 =" SEVERITY note;
		a_in <= O"4";
		b_in <= O"2";
		c_in <= '0';
		WAIT FOR stimulus_step_c;
		led7seg_show_big(an_out, seg_out);

		REPORT "7 + 7 + 1 =" SEVERITY note;
		a_in <= O"7";
		b_in <= O"7";
		c_in <= '1';
		WAIT FOR stimulus_step_c;
		led7seg_show_big(an_out, seg_out);

		-- Testujeme Adder3
		REPORT "Testing Adder3..." SEVERITY note;
		FOR a IN 0 TO 7 LOOP
			FOR b IN 0 TO 7 LOOP
				FOR c IN 0 TO 1 LOOP
					a_in <= std_logic_vector(to_unsigned(a, 3));
					b_in <= std_logic_vector(to_unsigned(b, 3));
					c_in <= std_logic(to_unsigned(c, 1)(0));
					WAIT FOR stimulus_step_c;

					--led7seg_show(an_out, seg_out);
					ASSERT(dut_sum_result = std_logic_vector(to_unsigned(a + b + c, 4)))
					 REPORT to_string(a) & "+" & to_string(b) & "+" & to_string(c) & " = " &
					  to_string(to_integer(unsigned(dut_sum_result))) SEVERITY error;
				END LOOP;
			END LOOP;
		END LOOP;

		-- Vynulujeme vstupy
		a_in <= (OTHERS => '0');
		b_in <= (OTHERS => '0');
		c_in <= '0';
		WAIT FOR stimulus_step_c;

		REPORT "Test done." SEVERITY note;
		WAIT;
	END PROCESS;
END Behavioral;
